`timescale 10ns/1ns
module and_gate(
	input A,
  	input B,
  	output out
);
  
  and A1 (out, A, B);
  
endmodule